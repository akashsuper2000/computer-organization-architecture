// module hey;
// wire c;
// reg a,b;
// hello mygate(.a(a), .b(b), .c(c));
// initial
// begin

// $monitor("%b & %b = %b", a,b,c);
// a = 0;
// b = 0;
// #1
// a = 0;
// b = 1;
// #1
// a = 1;
// b = 0;
// #1
// a = 1;
// b = 1;

// end
// endmodule






// module hey;
// wire c,d;
// reg a,b,cin;
// hello mygate(.a(a), .b(b), .cin(cin), .c(c), .d(d));
// initial
// begin

// $monitor("%b & %b & %b = %b, %b", a,b,cin,c,d);
// a = 0;
// b = 0;
// cin = 0;
// #1
// a = 0;
// b = 1;
// cin = 0;
// #1
// a = 1;
// b = 0;
// cin = 0;
// #1
// a = 1;
// b = 1;
// cin = 0;
// #1
// a = 0;
// b = 0;
// cin = 1;
// #1
// a = 0;
// b = 1;
// cin = 1;
// #1
// a = 1;
// b = 0;
// cin = 1;
// #1
// a = 1;
// b = 1;
// cin = 1;

// end
// endmodule






// module hey;
// wire c,d;
// reg a,b;
// hello mygate(.a(a), .b(b), .c(c), .d(d));
// initial
// begin

// $monitor("%b & %b = %b %b", a,b,c,d);
// a = 0;
// b = 0;
// #1
// a = 0;
// b = 1;
// #1
// a = 1;
// b = 0;
// #1
// a = 1;
// b = 1;

// end
// endmodule







// module hey;
// wire c,d;
// reg a,b,cin;
// hello mygate(.a(a), .b(b), .cin(cin), .c(c), .d(d));
// initial
// begin

// $monitor("%b & %b & %b = %b, %b", a,b,cin,c,d);
// a = 0;
// b = 0;
// cin = 0;
// #1
// a = 0;
// b = 1;
// cin = 0;
// #1
// a = 1;
// b = 0;
// cin = 0;
// #1
// a = 1;
// b = 1;
// cin = 0;
// #1
// a = 0;
// b = 0;
// cin = 1;
// #1
// a = 0;
// b = 1;
// cin = 1;
// #1
// a = 1;
// b = 0;
// cin = 1;
// #1
// a = 1;
// b = 1;
// cin = 1;

// end
// endmodule