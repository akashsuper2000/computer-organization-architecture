// module hello(a,b,c,d); 	
// input a,b;
// output c,d;
// wire ca, cb, cc, cd;

// xor(c,a,b);
// and(d,a,b);

// endmodule



// module hello(a,b,cin,c,d); 	
// input a,b,cin;
// output c,d;
// wire ca, cb, cc, cd;

// xor(ca,a,b);
// and(cb,a,b);
// xor(c,cin,ca);
// and(cc,ca,cin);
// or(d,cb,cc);

// endmodule



// module hello(a,b,c,d); 	
// input a,b;
// output c,d;
// wire ca, cb, cc, cd;

// xor(c,a,b);
// not(ca,a);
// and(d,ca,b);

// endmodule



// module hello(a,b,cin,c,d); 	
// input a,b,cin;
// output c,d;
// wire ca, cb, cc, cd;

// xor(ca,a,b);
// and(cb,a,b);
// xor(c,cin,ca);
// and(cc,ca,cin);
// or(d,cb,cc);

// endmodule